module processor();

endmodule