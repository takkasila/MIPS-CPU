module controller (
	, output reg RegDst
	, output reg Branch
	, output reg MemRead
	, output reg MemtoReg
	, output reg MemWrite
	, output reg ALUSrc
	, output reg RegWrite
	, output reg [5:0] ALUSelect_out
	, input [5:0] OPCode_in
	, input [5:0] ALUSelect_in);

	

endmodule